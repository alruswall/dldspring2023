module gol(start, clk, outGrid)
 input start;
 output [63:0] outGrid;
datapath prog(currentGrid, nextGrid)































endmodule